// CONFIDENTIAL AND PROPRIETARY INFORMATION
// Copyright 1998-2012 ARC International (Unpublished)
// All Rights Reserved.
//
// This document, material and/or software contains confidential
// and proprietary information of ARC International and is
// protected by copyright, trade secret and other state, federal,
// and international laws, and may be embodied in patents issued
// or pending.  Its receipt or possession does not convey any
// rights to use, reproduce, disclose its contents, or to
// manufacture, or sell anything it may describe.  Reverse
// engineering is prohibited, and reproduction, disclosure or use
// without specific written authorization of ARC International is
// strictly forbidden.  ARC and the ARC logotype are trademarks of
// ARC International.
// 
// ARC Product:  ARC 600 Architecture v4.9.7
// File version:  600 Architecture IP Library version 4.9.7, file revision 
// ARC Chip ID:  0
//
// Description:
//
// This module contains all the necessary logic for all debug
// extensions in the ARC.
//  
//  This file contains the debug extensions for:
// 
// 
//  L indicates a latched signal and U indicates a signal produced by
//  logic.
//
//======================= Inputs to this block =======================--
// 
//  aux_access       U Auxiliary Access. This signal is flagged by the
//                   host to inform the ARC that the address supplied on
//                   h_addr[31:0] applies to the auxiliary register set. 
// 
//  aux_addr[31:0]   U Auxiliary Register Address. This is produced by 
//                   the hostif.v, from the host address when the ARC
//                   is halted (en = '0') or from source 1 from pipeline
//                   stage 3, when the ARC is running. Width of decode is
//                   set by AUXDECSZ in extutil.v. 
// 
//  aux_dataw[31:0]  U Auxiliary Write Data. The auxiliary register bus 
//                   write data value is latched into auxiliary register
//                   specified by aux_addr[31:0] at the end of the cycle
//                   when aux_write is true. This is generated by 
//                   hostif.v, either from the host's write data bus 
//                   when the ARC is halted (en = '0') or from source 1
//                   from pipeline stage 3, when the ARC is running.
// 
//  aux_read         U Auxiliary Read. This signal indicates that a read 
//                   is taking place on this cycle. This is initiated
//                   either by an LR instruction when the ARC is running,
//                   or by a host read when the ARC is halted (for single 
//                   access aux registers). The data stored at location
//                   aux_addr[31:0] should be placed on drx_reg[31:0].
//                   The xreg_hit signal should be asserted if the
//                   register in question is recognised as a valid
//                   extension auxiliary register. For dual access
//                   registers, aux_regs.v and hostif.v will select
//                   the correct data values to go to the ARC and the
//                   host.
// 
//  aux_write        U Auxiliary Write. This signal indicates that a
//                   write (either from the ARC or host) is being
//                   performed to the auxiliary register specified on 
//                   aux_addr[31:0] on this cycle. This signal is set by
//                   hostif.v by a SR instruction when the ARC is
//                   running or a host when it is halted. The data 
//                   supplied by aux_dataw[31:0] should be latched into
//                   register specified by aux_addr[31:0] at the end of
//                   the cycle. For dual access extension registers,
//                   writes are ignored from regular auxiliary register
//                   bus aux_write, aux_addr(), and aux_dataw() when the
//                   ARC is halted.
// 
//  currentpc_nxt    U Pre-latch PC value. This is the value of program
//                   counter which corresponds to the ifetch_aligned 
//                   signal. It is latched by the ARC onto currentpc_r,
//                   and used by the processor.
//
//  currentpc_r      This is the latched value of the pc which is
//                   currently being used by stage 1 to fetch the next
//                   instruction. 
// 
//  dwr[]            Data value to be stored to memory. It is latched
//                   stval from the ARC interface. The value is latched
//                   when en2='1', i.e. the pipeline is not stalled.
// 
//  en               L Global enable. This is true when the ARC is
//                   running in normal operation.
// 
//  en1              U Stage 2 pipeline latch control. True when an
//                   instruction is being latched into pipeline stage 2.
//                   This will be true at different times to pcen, as it
//                   allows junk instructions to be latched into the
//                   pipeline.
//                   *** A feature of this signal is that it will allow
//                   an instruction be clocked into stage 2 even when
//                   stage 3 is halted, provided that stage 2 contains
//                   a killed instruction (i.e. p2iv = '0'). This is
//                   called a 'catch-up'. ***
// 
//  en2              U Pipeline stage 2 enable. When this signal is true,
//                   the instruction in stage 2 can pass into stage 3 at
//                   the end of the cycle. When it is false, it will
//                   hold up stage 2 and stage 1 (pcen).
// 
//  en3              U Pipeline stage 3 enable. When this signal is true,
//                   the instruction in stage 3 can pass into stage 4 at
//                   the end of the cycle. When it is false, it will
//                   probably hold up stages one (pcen), two (en2), and
//                   three. It is set in the rctl.v block.
//                   
//  h_addr[31:0]     L Host Address. This is a longword-granularity
//                   address latched by the host before being presented
//                   to the register module. This is a 32-bit address (it
//                   may be smaller, but packed with zeroes) from the
//                   host which is used to access registers in the ARC in
//                   conjuction with aux_access and core_access. The
//                   width of the decode applied to this 32-bit quantity
//                   is defined by the AUXDECSZ constant, found in
//                   extutil.v. It is defined as being a 32-bit bus at
//                   this level to maintain compatibility with the LR and 
//                   SR instructions which can generate a 32-bit value
//                   for the address to be used for auxiliary register
//                   accesses.
// 
//  h_dataw[31:0]    L Host Write Data. This bus carries the data which
//                   is to be stored into registers in the ARC or core 
//                   extensions. It is latched by the host as is the
//                   address, h_addr[31:0].
//                   
//  h_read           U Host Read. When the host signals h_read is true, 
//                   this signal indicates that a host read is taking
//                   place, and the register module should latch the data
//                   on h_dataw[31:0] at the end of the cycle.
// 
//  h_write          U Host Write. When the host signals h_write is true, 
//                   this signal indicates that a host write is taking
//                   place, and the register module should latch the data
//                   on h_dataw[31:0] at the end of the cycle.
// 
//  ifetch           U This signal, similar to pcen, indicates to the
//                   memory controller that a new instruction is
//                   required, and should be fetched from memory from the
//                   address which will be clocked into currentpc_r[31:0]
//                   at the end of the cycle. It is also true for one
//                   cycle when the processor has been started following
//                   a reset, in order to get the ball rolling.
//                   An instruction fetch will also be issued if the host
//                   changes the program counter when the ARC is halted,
//                   provided it is not directly after a reset.
//                   The ifetch signal will never be set true whilst the
//                   memory controller is in the process of doing an
//                   instruction fetch, so it may be used by the memory
//                   controller as an acknowledgement of instruction
//                   receipt.
// 
//  ivalid_aligned   U Qualifying signal for p1iw[31:0]. When it is low,
//                   this indicates that the m/c has not been able to
//                   fetch the requested opcode, and that the program
//                   counter should not be incremented. The pipeline
//                   might be stalled, depending upon whether the
//                   instruction in stage 2 needs to look at the
//                   instruction in stage 1. When it is true, the
//                   instruction is clocked into pipeline stage 2
//                   provided that the pipeline is able to move on.
// 
//  ldvalid          U From LSU. This signal is set true by the LSU to
//                   indicate that a delayed load writeback WILL occur on
//                   the next cycle. If the instruction in stage 3 wishes
//                   to perform a writeback, then pipeline stage 1, 2 and
//                   3 will be held. If the instruction is stage 3 is
//                   invalid, or does not want to write a value into the
//                   core register set for some reason, then the
//                   instructions in stages 1 and 2 will move into 2 and
//                   3 respectively, and the instruction that was in
//                   stage 3 will be replaced in stage 4 by the delayed
//                   load writeback. 
//                   ** Note that delayed load writebacks WILL complete,
//                   even if the processor is halted (en=0). In this
//                   instance, the host may be held off for a cycle
//                   (hold_host) if it is attempting to access the core
//                   registers. **
// 
//  mc_addr[]        The result of the adder unit. Goes to LSU, to be 
//                   latched by the memory controller.
// 
//  mstore           U This signal indicates to the LSU that there is a
//                   valid store instruction in stage 3.
// 
//  p2limm           U From rctl.v. This is used by the actionpoint
//                   debugging system when selected to qualify the value
//                   of the PC at stage one of the pipeline. The limm
//                   data is considered to be at the same the value
//                   address as the instruction it is associated with
//                   with regards to the debugger.
// 
//  p2opcode         L Opcode word. This bus contains the instruction
//                   word which is being executed by stage 2. It must be
//                   qualified by p2iv.
// 
//  p2iv             L Opcode valid. This signal is used to indicate that 
//                   the opcode in pipeline stage 2 is a valid
//                   instruction. The instruction may not be valid if a
//                   junk instruction has been allowed to come into the
//                   pipeline in order to allow the pipeline to continue
//                   running when an instruction cannot be fetched by the
//                   memory controller.
// 
//  kill_p1_a     U This signal indicates that the delay slot
//                   mechanism of the jump instruction currently in stage 
//                   2 is requesting that the next instruction be killed
//                   before it gets into stage 2. This signal is produced 
//                   from a decode for a jump instruction code, the 
//                   condition-true signal, p2iv and the delay-slot field
//                   in the instruction. This signal relies on the delay
//                   slot instruction being present in stage 1 before
//                   stage 2 can move on. This is handled elsewhere by
//                   this file.
// 
//  kill_p2_a        Kill Stage 2. This is asserted true when the
//                   instructin in stage 2 should be killed.
//
//  wba[5:0]         L This bus carries the address of the register to
//                   which the data on wbdata[31:0] is to be written at
//                   the end of the cycle if wben is true. It is produced
//                   during stage 3 and takes account of delayed load
//                   register writeback (taking a value from the LSU), 
//                   LD/ST address writeback (address from the B or C 
//                   field), and normal ALU operation destination
//                   addresses (instruction A field).
// 
//  wbdata[31:0]     L This is the bus which carries the latched (stage
//                   4) data to be written into the register file. This
//                   result is selected from numerous ALU results,
//                   delayed load register writebacks, and LR results.
//                   It is written into the register file at the end of
//                   the cycle if wben is true.
// 
//  wben             L This signal is the enable signal which determines
//                   whether the data on wbdata[31:0] is written into the 
//                   register file at stage 4. It is produced in stage 3
//                   and takes into account delayed load writebacks, 
//                   cancelled instructions, and instructions which are
//                   not to be executed due to the cc result being false,
//                   amongst other things.
// 
//======================== Output from this block ====================--
// 
//  actionpt_pc_addr_r
//                   L Actionpoint PC Address.
//
//  actionpt_status_r
//                   L Actionpoint Value. This registered bus can be
//                   read by the debugger from within the debug register 
//                   when the ARC has been halted by an actionpoint to 
//                   determine which one was responsible. There is a bit
//                   for each actionpoint in the system.
// 
//  actionpt_hit_a   U Actionpoint Valid. This signals to the ARC that it
//                   should be halted since a valid actionpoint has been
//                   set when it is true.
// 
//  en_debug_r       This flag is the Enable Debug flag (ED), bit 24 in
//                   the DEBUG register. It enables the debug extensions
//                   when it is set. When it is cleared the debug
//                   extensions are switched off by gating the debug
//                   clock, but only if the option clock gating has been
//                   selected.
//
//====================================================================--
//

module debug_exts (clk,
                   clk_debug,
                   clk_ungated,
                   rst_a,                   
                   ivic,                   
                   p2b_iv,
                   p2_iw_r,
                   actionpt_pc_brk_a,
                   p2_brcc_instr_a,
                   p3_brcc_instr_a,
                   p2_ap_stall_a,
                   p2b_jmp_holdup_a,
                   en,
                   aux_access,
                   aux_read,
                   aux_write,
                   core_access,
                   h_addr,
                   h_dataw,
                   h_write,
                   h_read,
                   en1,
                   en2,
                   en2b,
                   en3,
                   ivalid_aligned,
                   mload2b,
                   mstore2b,
                   mwait,
                   p2limm,
                   p2iv,
                   p2opcode,
                   p2subopcode,
                   currentpc_r,
                   p1iw,
                   mc_addr,
                   dwr,
                   drd,
                   aux_addr,
                   aux_dataw,
                   aux_datar,
                   ap_param0,
                   ap_param1,
                   ivalid,
                   kill_tagged_p1,
                   kill_p2_a,
                   mload,
                   mstore,
                   ldvalid,
                   ap_param0_read,
                   ap_param0_write,
                   ap_param1_read,
                   ap_param1_write,
// <add more signals as appropriate>

//Signals required for extensions are inserted here. The automatic
//hierarchy generation system can be used to create the structural
//HDL to tie all the components together, provided that certain
//naming and usage rules are followed. Please see the document
//'Automatic Hierarchy Generator' - $ARCHOME/arc/docs/hiergen.pdf
//

                   actionhalt,
                   actionpt_status_r,
                   ap_ahv0,
                   ap_ahv1,
                   ap_ahv2,
                   ap_ahv3,
                   ap_ahv4,
                   ap_ahv5,
                   ap_ahv6,
                   ap_ahv7,
                   ap_ahc0,
                   ap_ahc1,
                   ap_ahc2,
                   ap_ahc3,
                   ap_ahc4,
                   ap_ahc5,
                   ap_ahc6,
                   ap_ahc7,
                   ap_ahm0,
                   ap_ahm1,
                   ap_ahm2,
                   ap_ahm3,
                   ap_ahm4,
                   ap_ahm5,
                   ap_ahm6,
                   ap_ahm7,
                   actionpt_hit_a,
                   actionpt_swi_a,
                   en_debug_r);

`include "arcutil_pkg_defines.v"
`include "arcutil.v"
`include "extutil.v"
`include "xdefs.v"

//Extra include files required for extensions are inserted here.

input   clk;        // core clock
input   clk_ungated; // ungated core clock
input   clk_debug;  // debug clock
input   rst_a;      // system reset 
input   en;         // system go

// Debugger Access via Host Interface
// 
input   aux_access; 
input   aux_read; 
input   aux_write; 
input   core_access; 
input   [31:0] h_addr; 
input   [31:0] h_dataw; 
input   h_write; 
input   h_read;

input   ivic; 
input   en1; 
input   en2; 
input   en2b; 
input   en3; 
input   ivalid_aligned; 
input   mload2b; 
input   mstore2b; 
input   mwait; 
input   p2limm; 
input   p2iv; 
input   [4:0] p2opcode;
input   [5:0] p2subopcode;

// Actionpoint Data Sources
// 
input   [PC_MSB:0] currentpc_r; 
input   [31:0] p1iw;
input   [31:0] mc_addr; 
input   [31:0] dwr; 
input   [31:0] drd; 
input   [31:0] aux_addr; 
input   [31:0] aux_dataw; 
input   [31:0] aux_datar; 
input   [31:0] ap_param0;
input   [31:0] ap_param1;

// Actionpoint Data Sources Qualifiers
// 
input   ivalid;
input   kill_tagged_p1;
input   kill_p2_a;
input   p2b_jmp_holdup_a;
input   mload; 
input   mstore; 
input   ldvalid; 
input   ap_param0_read;
input   ap_param0_write;
input   ap_param1_read;
input   ap_param1_write;
input   p2b_iv;
input   [INSTR_UBND:0] p2_iw_r;
input   p2_brcc_instr_a;
input   p3_brcc_instr_a;



// Actionpoint Debug Hardware signals
//
input   actionhalt;

output  [NUM_APS - 1:0] actionpt_status_r; 
output  [31:0] ap_ahv0;
output  [31:0] ap_ahv1;
output  [31:0] ap_ahv2;
output  [31:0] ap_ahv3;
output  [31:0] ap_ahv4;
output  [31:0] ap_ahv5;
output  [31:0] ap_ahv6;
output  [31:0] ap_ahv7;
output  [31:0] ap_ahc0;
output  [31:0] ap_ahc1;
output  [31:0] ap_ahc2;
output  [31:0] ap_ahc3;
output  [31:0] ap_ahc4;
output  [31:0] ap_ahc5;
output  [31:0] ap_ahc6;
output  [31:0] ap_ahc7;
output  [31:0] ap_ahm0;
output  [31:0] ap_ahm1;
output  [31:0] ap_ahm2;
output  [31:0] ap_ahm3;
output  [31:0] ap_ahm4;
output  [31:0] ap_ahm5;
output  [31:0] ap_ahm6;
output  [31:0] ap_ahm7;
output  p2_ap_stall_a;
output  actionpt_pc_brk_a;
output  actionpt_hit_a; 
output  actionpt_swi_a; 
output  en_debug_r;


wire    [NUM_APS - 1:0] actionpt_status_r; 
wire    actionpt_hit_a;
wire    en_debug_r;
wire    i_actionpt_hit_a;
wire    i_actionpt_swi_a;

// Signal declarations for extensions to be added.

// ====================== Debug Modes Inserted Here ===================--
// 
// Drive this signal (to debug.v) when the actionpoint extension is
// not selected.


//Drive this signal (to flags.v) when the actionpoint extension is
//not selected.
//
assign actionpt_hit_a      = i_actionpt_hit_a;
assign actionpt_swi_a      = i_actionpt_swi_a;

// Debug extension logic functions are inserted here.

// ==================== Components Instantiated Below =================--
// 
// Debug component instantiations are inserted here.
   actionpoints U_actionpoints (
   .clk_ungated(clk_ungated), 
   .clk_debug(clk_debug), 
   .rst_a(rst_a), 
   .en(en),
   .kill_p2_a(kill_p2_a),
   .en1(en1),
   .en2(en2),
   .ivic(ivic),
   .actionpt_pc_brk_a(actionpt_pc_brk_a),
   .p2_brcc_instr_a(p2_brcc_instr_a),
   .p3_brcc_instr_a(p3_brcc_instr_a),
   .p2_ap_stall_a(p2_ap_stall_a),
   .p2b_jmp_holdup_a(p2b_jmp_holdup_a),       
   .p2_iw_r(p2_iw_r), 
   .currentpc_r(currentpc_r), 
   .mc_addr(mc_addr), 
   .dwr(dwr), 
   .drd(drd), 
   .aux_addr(aux_addr), 
   .aux_dataw(aux_dataw), 
   .aux_datar(aux_datar),
   .h_addr(h_addr),
   .h_dataw(h_dataw),
   .h_write(h_write ),
   .ap_param0(ap_param0), 
   .ap_param1(ap_param1), 
   .p2iv(p2iv),
   .p2b_iv(p2b_iv), 
   .mload(mload), 
   .mstore(mstore), 
   .ldvalid(ldvalid), 
   .aux_write(aux_write),
   .aux_read(aux_read), 
   .ap_param0_read(ap_param0_read), 
   .ap_param0_write(ap_param0_write), 
   .ap_param1_read(ap_param1_read), 
   .ap_param1_write(ap_param1_write), 
   .aux_access(aux_access),
   .actionhalt(actionhalt),
   .ap_ahv0(ap_ahv0), 
   .ap_ahv1(ap_ahv1), 
   .ap_ahv2(ap_ahv2), 
   .ap_ahv3(ap_ahv3), 
   .ap_ahv4(ap_ahv4), 
   .ap_ahv5(ap_ahv5), 
   .ap_ahv6(ap_ahv6), 
   .ap_ahv7(ap_ahv7), 
   .ap_ahc0(ap_ahc0),
   .ap_ahc1(ap_ahc1),
   .ap_ahc2(ap_ahc2),
   .ap_ahc3(ap_ahc3),
   .ap_ahc4(ap_ahc4),
   .ap_ahc5(ap_ahc5),
   .ap_ahc6(ap_ahc6),
   .ap_ahc7(ap_ahc7),
   .ap_ahm0(ap_ahm0),
   .ap_ahm1(ap_ahm1),
   .ap_ahm2(ap_ahm2),
   .ap_ahm3(ap_ahm3),
   .ap_ahm4(ap_ahm4),
   .ap_ahm5(ap_ahm5),
   .ap_ahm6(ap_ahm6),
   .ap_ahm7(ap_ahm7),
   .actionpt_status_r(actionpt_status_r), 
   .actionpt_swi_a(i_actionpt_swi_a), 
   .actionpt_brk_a(i_actionpt_hit_a), 
   .en_debug_r(en_debug_r)); 

endmodule // module debug_exts

