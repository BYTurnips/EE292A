// CONFIDENTIAL AND PROPRIETARY INFORMATION
// Copyright 1996-2012 ARC International (Unpublished)
// All Rights Reserved.
//
// This document, material and/or software contains confidential
// and proprietary information of ARC International and is
// protected by copyright, trade secret and other state, federal,
// and international laws, and may be embodied in patents issued
// or pending.  Its receipt or possession does not convey any
// rights to use, reproduce, disclose its contents, or to
// manufacture, or sell anything it may describe.  Reverse
// engineering is prohibited, and reproduction, disclosure or use
// without specific written authorization of ARC International is
// strictly forbidden.  ARC and the ARC logotype are trademarks of
// ARC International.
// 
// ARC Product:  ARC 600 Architecture v4.9.7
// File version:  600 Architecture IP Library version 4.9.7, file revision 
// ARC Chip ID:  0
//
// Description:
//
// This module contains all the necessary logic to control the interrupts
// in the ARC600.
// 
// The ARC600 interrupt system can be extended to provide altogether 29
// interrupt lines. There are still only two priority levels, level 1
// (low priority) and level 2 (medimum priority) but the interrupts
// priority levels of each interrupt signal is now programmable
// on-the-fly through an auxiliary register.
//  
// There is a relatively large number of interrupt signals that need to 
// go through a priority encoder to select the highest priority active 
// interrupt. A priority encoder with more than 24 lines can produce a
// critical path in the system. Thus the encoder is now pipelined in
// two stages. This adds to the number of flipflops in this module but
// ensures that no new critical path is introduced in the system. As a
// side effect, the detection of an interrupt has now an added one cycle
// latency.
// 
// ========================= Inputs to this block =====================--
// 
//    clk_ungated The core ungated clock signal.
// 
//    rst_a       The global system reset signal.
// 
//    aux_write   From auxiliary unit to indicate that a write to an
//                auxiliary register is happening. The logic in this 
//                module checks for the matching register address and if
//                so then allows the  update to the selected register to
//                take place.
// 
//   aux_addr     From auxiliary unit to carry the address of the aux reg
//                that is being accessed. The address is compared to the 
//                int_unit aux register addresses and if matched then the 
//                selected register is updated with the aux data value.
// 
//   aux_wdata    From the auxiliary unit that carries the data value for 
//                an aux register write. If the write strobe is asserted
//                and the aux address register matches one the addresses
//                in this unit then the int_unit aux register is updated
//                with the new data value on this bus.
// 
//    irq3        L Original low Priority (level 1) interrupt signals. 
//    irq4        These signals are level sensitive by default but can be
//    irq5        programmed to be pulse sensitive. The priority level
//                can also be programmed to be medium level.
// 
//    irq6        L Original med Priority (level 2) interrupt signals. 
//    irq7        These signals are level sensitive by default but can be
//                programmed to be pulse sensitive. The priority level
//                can also be programmed to be low level.
// 
//    irq8        L extension interrupt lines - level sensitive and low
//    ...         priority by default but can be programmed to be pulse 
//    irq31       sensitive or medium priority.
// 
//    instruction_error
//                Instruction error. Generated by rctl and handled as
//                an pulse-sensitive input in this file.
//                It comes from a decode of the instruction opcode field,
//                combined with the signal from the extensions which
//                indicates whether an extension instruction is valid or
//                not. It does not currently include a decode of the
//                instruction's C field for single-operand instructions.
// 
//    memory_error
//                U Memory error. pulse sensitive input for the memory 
//                controller to use.
// 
//    en1         U Stage 2 pipeline latch control. True when an
//                instruction is being latched into pipeline stage 2.
//                Will be true at different times to pcen, as it allows
//                junk instructions to be latched into the pipeline. Used
//                in this case to  allow the interrupt-flag/fantasy
//                instruction to be passed down the pipeline.
// 
//    en2         U Stage 3 pipeline latch control. Controls transition 
//                of instruction in stage 2 to stage 3. Used here for
//                passing the interrupt down the pipeline correctly.
// 
//    en3         U Stage 4 pipeline latch control. Controls transition
//                of instruction in stage 3 to stage 4. Used here for
//                passing the interrupt down the pipeline correctly.
// 
//    interrupt_holdoff
//                U Hold off interrupts during this cycle. This signal is
//                set true by rctl.v to prevent an interrupt-op from
//                being inserted when a jump is in stage 2 (no interrupts
//                during delay slots) or when an instruction which uses 
//                long immediate data is in stage 2. This signal (or a
//                similar one) will be used in pipectl to prevent junk
//                instructions being inserted into the pipeline when
//                there is an interdependancy between the instructions
//                in stage 2 and the instruction in stage 1. Note that
//                this signal includes p2iv.
// 
//    e1flag_r      L from flags.v. The level 1 interrupt mask bit. 
// 
//    e2flag_r      L from flags.v. The level 2 interrupt mask bit. 
// 
// ======================== Output from this block ====================--
//
//    p1int       U indicates that an interrupt has been detected, and an
//                interrupt-op will be inserted into stage 2 on the next
//                cycle, (subject to pipeline enables) setting p2int
//                true. This signal will have the effect of cancelling
//                the instruction currently being fetched by stage 1 by
//                causing p2iv to be set false at the end of the cycle
//                when p1int is true.
// 
//    p2int       L Indicates that an interrupt-op instruction is in
//                stage 2. This signal is used in coreregs.v to control
//                the placing of the pc onto a source bus for writing
//                back to the interrupt link registers, and by aux_regs
//                to insert the interrupt vector int_vec[] into the
//                program counter.
// 
//    p2ilev1     L Indicates that the interrupt-op instruction in stage
//                2 was caused by a level 1 interrupt (irq3,4,5). It is
//                used by the load/store unit to stall an interrupt at
//                stage 2 if any loads are pending to ilink1 or ilink2.
// 
//    p2bint      L Indicates that an interrupt-op instruction is in
//                stage 2B. 
// 
//    p2bilev1    L Indicates that the interrupt-op instruction in stage
//                2B was caused by a level 1 interrupt (irq3,4,5). 
// 
//    p3int       L Indicates that an interrupt-op instruction is in 
//                stage 3. This signal is used by flags.v, along with
//                the p3ilev1 signal to clear one or both of the
//                interrupt mask bits in the status register.
// 
//    p3ilev1     L Indicates that the interrupt-op instruction in stage
//                3 was caused by a level 1 interrupt (irq3,4,5) and that 
//                only the e1 bit should be cleared. When this signal is
//                not true when p3int is true, both e1 and e2 bits are 
//                cleared. Also used to supply the correct register
//                address for the link register writeback.
// 
//    p123int     U Indicates that there is an interrupt in stage 1,2 or
//                3. This signal is used by the clock generation module.
//                If the option clock gating was not chosen this signal
//                is removed during synthesis.
// 
//    aux_lev     To auxliary unit to indicate the current value of the
//                interrupt level priority for all the interrupts. The 
//                programmer can set the priority of low priority by
//                writing to an aux register which is decoded and 
//                processed in this unit.
// 
//    int_vec     U This is the interrupt vector supplied to the 
//                program counter. Each interrupt line has a different
//                vector associated with it. It is latched into the PC
//                at the end of the cycle when p2int is true.
// 
//====================================================================--
//
module int_unit (clk_ungated,
                 rst_a,
                 irq,
                 instruction_error,
                 int_vector_base_r,
                 memory_error,
                 misaligned_int,
                 en1,
                 en2,
                 en2b,
                 en3,
                 interrupt_holdoff,
                 flagu_block,
                 e1flag_r,
                 e2flag_r,
                 aux_access,
                 aux_addr,
                 aux_dataw,
                 aux_write,
                 h_write,
                 h_addr,
                 h_dataw,
		 hold_int_st2_a,

                 int_vec,
                 p1int,
                 p2int,
                 p2bint,
                 p2ilev1,
                 p2bilev1,
                 p3int,
                 p3ilev1,
                 p123int,
                 aux_lv12,
                 aux_hint,
                 aux_lev);

`include "arcutil_pkg_defines.v" 
`include "arcutil.v" 
`include "extutil.v" 
`include "xdefs.v" 

input                       clk_ungated; 
input                       rst_a; 
input   [31:3]              irq; 
input                       instruction_error; 
input   [PC_MSB : `INT_BASE_LSB] int_vector_base_r; 
input                       memory_error; 
input                       misaligned_int;
input                       en1; 
input                       en2; 
input                       en2b; 
input                       en3; 
input                       interrupt_holdoff; 
input                       flagu_block; 
input                       e1flag_r; 
input                       e2flag_r; 
input                       aux_access; 
input   [31:0]              aux_addr; 
input   [31:0]              aux_dataw; 
input                       aux_write; 
input                       h_write; 
input   [31:0]              h_addr; 
input   [31:0]              h_dataw; 
input                       hold_int_st2_a;

output  [PC_MSB:0]          int_vec; 
output                      p1int; 
output                      p2int; 
output                      p2bint; 
output                      p2ilev1; 
output                      p2bilev1; 
output                      p3int; 
output                      p3ilev1; 
output                      p123int; 
output  [1:0]               aux_lv12; 
output  [4:0]               aux_hint; 
output   [31:3] aux_lev; 
wire    [PC_MSB:0]          int_vec; 
wire                        p1int; 
wire                        p2int; 
wire                        p2bint; 
wire                        p2ilev1; 
wire                        p2bilev1; 
wire                        p3int; 
wire                        p3ilev1; 
wire                        p123int; 
wire    [1:0]               aux_lv12; 
wire    [4:0]               aux_hint; 
wire    [31:3] aux_lev; 
reg [28:0]   i_swi_cancel_a;

//  INT_UNIT ARCHITECTURE
//
//  interrupt state constants
//
parameter S_IRQ0 = 5'b 00000; //  s_idle
parameter S_IRQ1 = 5'b 00001; //  s_mem
parameter S_IRQ2 = 5'b 00010; //  s_ins
parameter S_IRQ3 = 5'b 00011; 
parameter S_IRQ4 = 5'b 00100; 
parameter S_IRQ5 = 5'b 00101; 
parameter S_IRQ6 = 5'b 00110; 
parameter S_IRQ7 = 5'b 00111; 
parameter S_IRQ8 = 5'b 01000; 
parameter S_IRQ9 = 5'b 01001; 
parameter S_IRQ10 = 5'b 01010; 
parameter S_IRQ11 = 5'b 01011; 
parameter S_IRQ12 = 5'b 01100; 
parameter S_IRQ13 = 5'b 01101; 
parameter S_IRQ14 = 5'b 01110; 
parameter S_IRQ15 = 5'b 01111; 

parameter S_IRQ16 = 5'b 10000; 
parameter S_IRQ17 = 5'b 10001; 
parameter S_IRQ18 = 5'b 10010; 
parameter S_IRQ19 = 5'b 10011; 
parameter S_IRQ20 = 5'b 10100; 
parameter S_IRQ21 = 5'b 10101; 
parameter S_IRQ22 = 5'b 10110; 
parameter S_IRQ23 = 5'b 10111; 
parameter S_IRQ24 = 5'b 11000; 
parameter S_IRQ25 = 5'b 11001; 
parameter S_IRQ26 = 5'b 11010; 
parameter S_IRQ27 = 5'b 11011; 
parameter S_IRQ28 = 5'b 11100; 
parameter S_IRQ29 = 5'b 11101; 
parameter S_IRQ30 = 5'b 11110; 
parameter S_IRQ31 = 5'b 11111; 

//  Internal signals
//
//  Auxiliary registers
//
reg     [`INT_BASE_LSB_1:0] i_int_vec_a; 

reg     [31:3] i_aux_lev_r; 

//  Sticky flag that is set in hardware to indicate if a level 1
//  interrupt is taken. The flag should be reset in software.
//
reg     [1:0] i_aux_lev12_r; 

//  Five bits to encode the software triggered interrupt
//
reg     [4:0] i_aux_hint_r; 

//  Auxiliary lines for software driven interrupts
//
reg    [31:3] i_aux_hint_a; 

//  interrupt signals and registers
//
wire    [31:1] i_irq_a; 

reg     i_irq1_r; 
reg     i_irq2_r; 
reg     i_irq3_r; 
reg     i_irq4_r; 
reg     i_irq5_r; 
reg     i_irq6_r; 
reg     i_irq7_r; 
reg     i_irq8_r; 
reg     i_irq9_r; 
reg     i_irq10_r; 
reg     i_irq11_r; 
reg     i_irq12_r; 
reg     i_irq13_r; 
reg     i_irq14_r; 
reg     i_irq15_r; 

reg     i_irq16_r; 
reg     i_irq17_r; 
reg     i_irq18_r; 
reg     i_irq19_r; 
reg     i_irq20_r; 
reg     i_irq21_r; 
reg     i_irq22_r; 
reg     i_irq23_r; 
reg     i_irq24_r; 
reg     i_irq25_r; 
reg     i_irq26_r; 
reg     i_irq27_r; 
reg     i_irq28_r; 
reg     i_irq29_r; 
reg     i_irq30_r; 
reg     i_irq31_r; 

// Intermediate irq signals and states for stage 0,1 and 2
//
wire    [4:0] i_p0state0_nxt; 
wire    [4:0] i_p0state1_nxt; 
wire    [4:0] i_p0state2_nxt; 
wire    [4:0] i_p0state3_nxt; 
reg     [4:0] i_p0state0_r; 
reg     [4:0] i_p0state1_r; 
reg     [4:0] i_p0state2_r; 
reg     [4:0] i_p0state3_r; 
wire    [4:0] i_p1state_a; 
reg     [4:0] i_p2state_r; 

// Miscellanous internal signals
//
wire    i_blockout_a; 
wire    i_p1int_a; 
reg     i_p2bilevel1_r; 
wire    i_p2bint_nxt; 
reg     i_p2bint_r; 
wire    i_p2int_nxt; 
reg     i_p2int_r; 
reg     i_p2ilevel1_r; 
wire    i_p3int_nxt; 
reg     i_p3int_r; 
reg     i_p3ilevel1_r; 




// Select host interrupt
//
always @(
         i_aux_hint_r
         )
   begin : aux_hint_async_PROC
      case(i_aux_hint_r) 
        5'b 00011 : i_aux_hint_a = TWENTYNINE_ONE        ;
        5'b 00100 : i_aux_hint_a = TWENTYNINE_TWO        ;
        5'b 00101 : i_aux_hint_a = TWENTYNINE_THREE      ;
        5'b 00110 : i_aux_hint_a = TWENTYNINE_FOUR       ;
        5'b 00111 : i_aux_hint_a = TWENTYNINE_FIVE       ; 
        5'b 01000 : i_aux_hint_a = TWENTYNINE_SIX        ; 
        5'b 01001 : i_aux_hint_a = TWENTYNINE_SEVEN      ; 
        5'b 01010 : i_aux_hint_a = TWENTYNINE_EIGHT      ; 
        5'b 01011 : i_aux_hint_a = TWENTYNINE_NINE       ;
        5'b 01100 : i_aux_hint_a = TWENTYNINE_TEN        ;
        5'b 01101 : i_aux_hint_a = TWENTYNINE_ELEVEN     ;
        5'b 01110 : i_aux_hint_a = TWENTYNINE_TWELVE     ;
        5'b 01111 : i_aux_hint_a = TWENTYNINE_THIRTEEN   ;
        5'b 10000 : i_aux_hint_a = TWENTYNINE_FOURTEEN   ;
        5'b 10001 : i_aux_hint_a = TWENTYNINE_FIFTEEN    ;
        5'b 10010 : i_aux_hint_a = TWENTYNINE_SIXTEEN    ;
        5'b 10011 : i_aux_hint_a = TWENTYNINE_SEVENTEEN  ;
        5'b 10100 : i_aux_hint_a = TWENTYNINE_EIGHTEEN   ; 
        5'b 10101 : i_aux_hint_a = TWENTYNINE_NINETEEN   ; 
        5'b 10110 : i_aux_hint_a = TWENTYNINE_TWENTY     ; 
        5'b 10111 : i_aux_hint_a = TWENTYNINE_TWENTYONE  ; 
        5'b 11000 : i_aux_hint_a = TWENTYNINE_TWENTYTWO  ;
        5'b 11001 : i_aux_hint_a = TWENTYNINE_TWENTYTHREE;
        5'b 11010 : i_aux_hint_a = TWENTYNINE_TWENTYFOUR ;
        5'b 11011 : i_aux_hint_a = TWENTYNINE_TWENTYFIVE ;
        5'b 11100 : i_aux_hint_a = TWENTYNINE_TWENTYSIX  ;
        5'b 11101 : i_aux_hint_a = TWENTYNINE_TWENTYSEVEN;
        5'b 11110 : i_aux_hint_a = TWENTYNINE_TWENTYEIGHT;
        5'b 11111 : i_aux_hint_a = TWENTYNINE_TWENTYNINE ;  
        default   : i_aux_hint_a = THENTYNINE_ZERO       ;      
      endcase // case(l_aux_hit)
   end // block: i_aux_hit_mux
   

// An intermediate signal is created here which is true when:
//
//  a. The incoming interrupt signal is true
//
//  b. The intermediate signal was true on the last cycle.
//
// The intermediate signal is held low when the interrupt to 
// which it relates has been issued - i.e. has made it to stage 
// 2 of the pipeline. At this point blockout is asserted, so no 
// additional interrupts could be issued.
//
// Since the intermediate signal was held low on the previous 
// cycle, it will remain low until another pulse is received on 
// the incoming interrupt line.
//
// i_irq_a(0) is the reset exception and is handled differently.
//
assign i_irq_a[1] = ((memory_error | misaligned_int |
                    i_irq1_r) == 1'b 1 ) &
                  ( i_p2state_r != S_IRQ1 ) ? 1'b 1 : 
       1'b 0;

assign i_irq_a[2] = ( (instruction_error | i_irq2_r) == 1'b 1 ) &
                  ( i_p2state_r != S_IRQ2 ) ? 1'b 1 : 
       1'b 0;

assign i_irq_a[3] = ( (irq[3] | i_irq3_r | i_aux_hint_a[3]) == 1'b 1 ) & 
                  ( i_p2state_r != S_IRQ3 ) ? 1'b 1 : 
       1'b 0;

assign i_irq_a[4] = ( (irq[4] | i_irq4_r | i_aux_hint_a[4]) == 1'b 1 ) & 
                   ( i_p2state_r != S_IRQ4 ) ? 1'b 1 : 
       1'b 0;

assign i_irq_a[5] = ( (irq[5]  | i_irq5_r | i_aux_hint_a[5]) == 1'b 1 ) & 
                  ( i_p2state_r != S_IRQ5 ) ? 1'b 1 : 
       1'b 0;

assign i_irq_a[6] = ( (irq[6]  | i_irq6_r | i_aux_hint_a[6]) == 1'b 1 ) & 
                  ( i_p2state_r != S_IRQ6 ) ? 1'b 1 : 
       1'b 0;

assign i_irq_a[7] = ( (irq[7]  | i_irq7_r | i_aux_hint_a[7]) == 1'b 1 ) & 
                  ( i_p2state_r != S_IRQ7 ) ? 1'b 1 : 
       1'b 0;

assign i_irq_a[8] = ( (irq[8] | i_irq8_r | i_aux_hint_a[8]) == 1'b 1 ) & 
                   ( i_p2state_r != S_IRQ8 ) ? 1'b 1 : 
       1'b 0;
 
assign i_irq_a[9] = ( (irq[9] | i_irq9_r | i_aux_hint_a[9]) == 1'b 1 ) & 
                   ( i_p2state_r != S_IRQ9 ) ? 1'b 1 : 
       1'b 0;

assign i_irq_a[10] = ( (irq[10] | i_irq10_r | i_aux_hint_a[10]) == 1'b 1 ) & 
                   ( i_p2state_r != S_IRQ10 ) ? 1'b 1 : 
       1'b 0;

assign i_irq_a[11] = ( (irq[11] | i_irq11_r | i_aux_hint_a[11]) == 1'b 1 ) & 
                   ( i_p2state_r != S_IRQ11 ) ? 1'b 1 : 
       1'b 0;

assign i_irq_a[12] = ( (irq[12] | i_irq12_r | i_aux_hint_a[12]) == 1'b 1 ) & 
                   ( i_p2state_r != S_IRQ12 ) ? 1'b 1 : 
       1'b 0;

assign i_irq_a[13] = ( (irq[13] | i_irq13_r | i_aux_hint_a[13]) == 1'b 1 ) & 
                   ( i_p2state_r != S_IRQ13 ) ? 1'b 1 : 
       1'b 0;

assign i_irq_a[14] = ( (irq[14] | i_irq14_r | i_aux_hint_a[14]) == 1'b 1 ) & 
                   ( i_p2state_r != S_IRQ14 ) ? 1'b 1 : 
       1'b 0;

assign i_irq_a[15] = ( (irq[15] | i_irq15_r | i_aux_hint_a[15]) == 1'b 1 ) & 
                   ( i_p2state_r != S_IRQ15 ) ? 1'b 1 : 
       1'b 0;

assign i_irq_a[16] = (((irq[16] | i_irq16_r | i_aux_hint_a[16]) == 1'b 1) & 
                   (i_p2state_r != S_IRQ16)) ? 1'b 1 : 
       1'b 0;
assign i_irq_a[17] = (((irq[17] | i_irq17_r | i_aux_hint_a[17]) == 1'b 1) & 
                   (i_p2state_r != S_IRQ17)) ? 1'b 1 : 
       1'b 0;
assign i_irq_a[18] = (((irq[18] | i_irq18_r | i_aux_hint_a[18]) == 1'b 1) & 
                   (i_p2state_r != S_IRQ18)) ? 1'b 1 : 
       1'b 0;
assign i_irq_a[19] = (((irq[19] | i_irq19_r | i_aux_hint_a[19]) == 1'b 1) & 
                   (i_p2state_r != S_IRQ19)) ? 1'b 1 : 
       1'b 0;
assign i_irq_a[20] = (((irq[20] | i_irq20_r | i_aux_hint_a[20]) == 1'b 1) & 
                   (i_p2state_r != S_IRQ20)) ? 1'b 1 : 
       1'b 0;
assign i_irq_a[21] = (((irq[21] | i_irq21_r | i_aux_hint_a[21]) == 1'b 1) & 
                   (i_p2state_r != S_IRQ21)) ? 1'b 1 : 
       1'b 0;
assign i_irq_a[22] = (((irq[22] | i_irq22_r | i_aux_hint_a[22]) == 1'b 1) & 
                   (i_p2state_r != S_IRQ22)) ? 1'b 1 : 
       1'b 0;
assign i_irq_a[23] = (((irq[23] | i_irq23_r | i_aux_hint_a[23]) == 1'b 1) & 
                   (i_p2state_r != S_IRQ23)) ? 1'b 1 : 
       1'b 0;
assign i_irq_a[24] = (((irq[24] | i_irq24_r | i_aux_hint_a[24]) == 1'b 1) & 
                   (i_p2state_r != S_IRQ24)) ? 1'b 1 : 
       1'b 0;
assign i_irq_a[25] = (((irq[25] | i_irq25_r | i_aux_hint_a[25]) == 1'b 1) & 
                   (i_p2state_r != S_IRQ25)) ? 1'b 1 : 
       1'b 0;
assign i_irq_a[26] = (((irq[26] | i_irq26_r | i_aux_hint_a[26]) == 1'b 1) & 
                   (i_p2state_r != S_IRQ26)) ? 1'b 1 : 
       1'b 0;
assign i_irq_a[27] = (((irq[27] | i_irq27_r | i_aux_hint_a[27]) == 1'b 1) & 
                   (i_p2state_r != S_IRQ27)) ? 1'b 1 : 
       1'b 0;
assign i_irq_a[28] = (((irq[28] | i_irq28_r | i_aux_hint_a[28]) == 1'b 1) & 
                   (i_p2state_r != S_IRQ28)) ? 1'b 1 : 
       1'b 0;
assign i_irq_a[29] = (((irq[29] | i_irq29_r | i_aux_hint_a[29]) == 1'b 1) & 
                   (i_p2state_r != S_IRQ29)) ? 1'b 1 : 
       1'b 0;
assign i_irq_a[30] = (((irq[30] | i_irq30_r | i_aux_hint_a[30]) == 1'b 1) & 
                   (i_p2state_r != S_IRQ30)) ? 1'b 1 : 
       1'b 0;
assign i_irq_a[31] = (((irq[31] | i_irq31_r | i_aux_hint_a[31]) == 1'b 1) & 
                   (i_p2state_r != S_IRQ31)) ? 1'b 1 : 
       1'b 0;

// Process to register pulse sensitive interrupts and store the
// auxiliary write values coding: '0' = level , '1' = pulse
//
always @(posedge clk_ungated or posedge rst_a)
   begin : reg_irqs_PROC

   if (rst_a == 1'b 1)
      begin

   //  Reset stored intermediate signals & auxiliary registers
   //
      i_aux_lev_r <= 29'b00000000000000000000000011000;
      i_aux_hint_r <= 5'b 00000;    

   // The format of the logic for the interrupts represented below is
   // will cause synthesis tools to flag warnings. Note these can be
   // ignored since they appear when the interrupts are set to being
   // level sensitive.
   //
      if (MEM_IRQ_TYPE == IRQ_TYPE_LEVEL)
         begin
         i_irq1_r <= 1'b 0; 
         end
      if (INS_IRQ_TYPE == IRQ_TYPE_LEVEL)
         begin
         i_irq2_r <= 1'b 0; 
         end
      if (IRQ3_TYPE == IRQ_TYPE_LEVEL)
         begin
         i_irq3_r <= 1'b 0; 
         end
      if (IRQ4_TYPE == IRQ_TYPE_LEVEL)
         begin
         i_irq4_r <= 1'b 0; 
         end
      if (IRQ5_TYPE == IRQ_TYPE_LEVEL)
         begin
         i_irq5_r <= 1'b 0; 
         end
      if (IRQ6_TYPE == IRQ_TYPE_LEVEL)
         begin
         i_irq6_r <= 1'b 0; 
         end
      if (IRQ7_TYPE == IRQ_TYPE_LEVEL)
         begin
         i_irq7_r <= 1'b 0; 
         end
      if (IRQ8_TYPE == IRQ_TYPE_LEVEL)
         begin
         i_irq8_r <= 1'b 0; 
         end
      if (IRQ9_TYPE == IRQ_TYPE_LEVEL)
         begin
         i_irq9_r <= 1'b 0; 
         end
      if (IRQ10_TYPE == IRQ_TYPE_LEVEL)
         begin
         i_irq10_r <= 1'b 0;    
         end
      if (IRQ11_TYPE == IRQ_TYPE_LEVEL)
         begin
         i_irq11_r <= 1'b 0;    
         end
      if (IRQ12_TYPE == IRQ_TYPE_LEVEL)
         begin
         i_irq12_r <= 1'b 0;    
         end
      if (IRQ13_TYPE == IRQ_TYPE_LEVEL)
         begin
         i_irq13_r <= 1'b 0;    
         end
      if (IRQ14_TYPE == IRQ_TYPE_LEVEL)
         begin
         i_irq14_r <= 1'b 0;    
         end
      if (IRQ15_TYPE == IRQ_TYPE_LEVEL)
         begin
         i_irq15_r <= 1'b 0;    
         end

      if (IRQ16_TYPE == IRQ_TYPE_LEVEL) begin i_irq16_r <= 1'b 0;    end
      if (IRQ17_TYPE == IRQ_TYPE_LEVEL) begin i_irq17_r <= 1'b 0;    end
      if (IRQ18_TYPE == IRQ_TYPE_LEVEL) begin i_irq18_r <= 1'b 0;    end
      if (IRQ19_TYPE == IRQ_TYPE_LEVEL) begin i_irq19_r <= 1'b 0;    end
      if (IRQ20_TYPE == IRQ_TYPE_LEVEL) begin i_irq20_r <= 1'b 0;    end
      if (IRQ21_TYPE == IRQ_TYPE_LEVEL) begin i_irq21_r <= 1'b 0;    end
      if (IRQ22_TYPE == IRQ_TYPE_LEVEL) begin i_irq22_r <= 1'b 0;    end
      if (IRQ23_TYPE == IRQ_TYPE_LEVEL) begin i_irq23_r <= 1'b 0;    end
      if (IRQ24_TYPE == IRQ_TYPE_LEVEL) begin i_irq24_r <= 1'b 0;    end
      if (IRQ25_TYPE == IRQ_TYPE_LEVEL) begin i_irq25_r <= 1'b 0;    end
      if (IRQ26_TYPE == IRQ_TYPE_LEVEL) begin i_irq26_r <= 1'b 0;    end
      if (IRQ27_TYPE == IRQ_TYPE_LEVEL) begin i_irq27_r <= 1'b 0;    end
      if (IRQ28_TYPE == IRQ_TYPE_LEVEL) begin i_irq28_r <= 1'b 0;    end
      if (IRQ29_TYPE == IRQ_TYPE_LEVEL) begin i_irq29_r <= 1'b 0;    end
      if (IRQ30_TYPE == IRQ_TYPE_LEVEL) begin i_irq30_r <= 1'b 0;    end
      if (IRQ31_TYPE == IRQ_TYPE_LEVEL) begin i_irq31_r <= 1'b 0;    end

      if (MEM_IRQ_TYPE == IRQ_TYPE_PULSE)
         begin
         i_irq1_r <= 1'b 0; 
         end
      if (INS_IRQ_TYPE == IRQ_TYPE_PULSE)
         begin
         i_irq2_r <= 1'b 0; 
         end
      if (IRQ3_TYPE == IRQ_TYPE_PULSE)
         begin
         i_irq3_r <= 1'b 0; 
         end
      if (IRQ4_TYPE == IRQ_TYPE_PULSE)
         begin
         i_irq4_r <= 1'b 0; 
         end
      if (IRQ5_TYPE == IRQ_TYPE_PULSE)
         begin
         i_irq5_r <= 1'b 0; 
         end
      if (IRQ6_TYPE == IRQ_TYPE_PULSE)
         begin
         i_irq6_r <= 1'b 0; 
         end
      if (IRQ7_TYPE == IRQ_TYPE_PULSE)
         begin
         i_irq7_r <= 1'b 0; 
         end
      if (IRQ8_TYPE == IRQ_TYPE_PULSE)
         begin
         i_irq8_r <= 1'b 0; 
         end
      if (IRQ9_TYPE == IRQ_TYPE_PULSE)
         begin
         i_irq9_r <= 1'b 0; 
         end
      if (IRQ10_TYPE == IRQ_TYPE_PULSE)
         begin
         i_irq10_r <= 1'b 0;    
         end
      if (IRQ11_TYPE == IRQ_TYPE_PULSE)
         begin
         i_irq11_r <= 1'b 0;    
         end
      if (IRQ12_TYPE == IRQ_TYPE_PULSE)
         begin
         i_irq12_r <= 1'b 0;    
         end
      if (IRQ13_TYPE == IRQ_TYPE_PULSE)
         begin
         i_irq13_r <= 1'b 0;    
         end
      if (IRQ14_TYPE == IRQ_TYPE_PULSE)
         begin
         i_irq14_r <= 1'b 0;    
         end
      if (IRQ15_TYPE == IRQ_TYPE_PULSE)
         begin
         i_irq15_r <= 1'b 0;    
         end

      if (IRQ16_TYPE == IRQ_TYPE_PULSE) begin i_irq16_r <= 1'b 0;    end
      if (IRQ17_TYPE == IRQ_TYPE_PULSE) begin i_irq17_r <= 1'b 0;    end
      if (IRQ18_TYPE == IRQ_TYPE_PULSE) begin i_irq18_r <= 1'b 0;    end
      if (IRQ19_TYPE == IRQ_TYPE_PULSE) begin i_irq19_r <= 1'b 0;    end
      if (IRQ20_TYPE == IRQ_TYPE_PULSE) begin i_irq20_r <= 1'b 0;    end
      if (IRQ21_TYPE == IRQ_TYPE_PULSE) begin i_irq21_r <= 1'b 0;    end
      if (IRQ22_TYPE == IRQ_TYPE_PULSE) begin i_irq22_r <= 1'b 0;    end
      if (IRQ23_TYPE == IRQ_TYPE_PULSE) begin i_irq23_r <= 1'b 0;    end
      if (IRQ24_TYPE == IRQ_TYPE_PULSE) begin i_irq24_r <= 1'b 0;    end
      if (IRQ25_TYPE == IRQ_TYPE_PULSE) begin i_irq25_r <= 1'b 0;    end
      if (IRQ26_TYPE == IRQ_TYPE_PULSE) begin i_irq26_r <= 1'b 0;    end
      if (IRQ27_TYPE == IRQ_TYPE_PULSE) begin i_irq27_r <= 1'b 0;    end
      if (IRQ28_TYPE == IRQ_TYPE_PULSE) begin i_irq28_r <= 1'b 0;    end
      if (IRQ29_TYPE == IRQ_TYPE_PULSE) begin i_irq29_r <= 1'b 0;    end
      if (IRQ30_TYPE == IRQ_TYPE_PULSE) begin i_irq30_r <= 1'b 0;    end
      if (IRQ31_TYPE == IRQ_TYPE_PULSE) begin i_irq31_r <= 1'b 0;    end

      end

   else
      begin

      // Store last value of interrupt signal if pulse catching
      // is required. The value will be reset to zero when the
      // interrupt is issued, since the intermediate value
      // is held low when the correct interrupt is issued.
      //
      // i_irq_a (0) corresponds to reset exception.
      //
      if (MEM_IRQ_TYPE == IRQ_TYPE_LEVEL)
         begin
         i_irq1_r <= 1'b 0; 
         end
      if (INS_IRQ_TYPE == IRQ_TYPE_LEVEL)
         begin
         i_irq2_r <= 1'b 0; 
         end
      if (IRQ3_TYPE == IRQ_TYPE_LEVEL)
         begin
         i_irq3_r <= 1'b 0; 
         end
      if (IRQ4_TYPE == IRQ_TYPE_LEVEL)
         begin
         i_irq4_r <= 1'b 0; 
         end
      if (IRQ5_TYPE == IRQ_TYPE_LEVEL)
         begin
         i_irq5_r <= 1'b 0; 
         end
      if (IRQ6_TYPE == IRQ_TYPE_LEVEL)
         begin
         i_irq6_r <= 1'b 0; 
         end
      if (IRQ7_TYPE == IRQ_TYPE_LEVEL)
         begin
         i_irq7_r <= 1'b 0; 
         end
      if (IRQ8_TYPE == IRQ_TYPE_LEVEL)
         begin
         i_irq8_r <= 1'b 0; 
         end
      if (IRQ9_TYPE == IRQ_TYPE_LEVEL)
         begin
         i_irq9_r <= 1'b 0; 
         end
      if (IRQ10_TYPE == IRQ_TYPE_LEVEL)
         begin
         i_irq10_r <= 1'b 0;    
         end
      if (IRQ11_TYPE == IRQ_TYPE_LEVEL)
         begin
         i_irq11_r <= 1'b 0;    
         end
      if (IRQ12_TYPE == IRQ_TYPE_LEVEL)
         begin
         i_irq12_r <= 1'b 0;    
         end
      if (IRQ13_TYPE == IRQ_TYPE_LEVEL)
         begin
         i_irq13_r <= 1'b 0;    
         end
      if (IRQ14_TYPE == IRQ_TYPE_LEVEL)
         begin
         i_irq14_r <= 1'b 0;    
         end
      if (IRQ15_TYPE == IRQ_TYPE_LEVEL)
         begin
         i_irq15_r <= 1'b 0;    
         end

      if (IRQ16_TYPE == IRQ_TYPE_LEVEL) begin i_irq16_r <= 1'b 0;    end
      if (IRQ17_TYPE == IRQ_TYPE_LEVEL) begin i_irq17_r <= 1'b 0;    end
      if (IRQ18_TYPE == IRQ_TYPE_LEVEL) begin i_irq18_r <= 1'b 0;    end
      if (IRQ19_TYPE == IRQ_TYPE_LEVEL) begin i_irq19_r <= 1'b 0;    end
      if (IRQ20_TYPE == IRQ_TYPE_LEVEL) begin i_irq20_r <= 1'b 0;    end
      if (IRQ21_TYPE == IRQ_TYPE_LEVEL) begin i_irq21_r <= 1'b 0;    end
      if (IRQ22_TYPE == IRQ_TYPE_LEVEL) begin i_irq22_r <= 1'b 0;    end
      if (IRQ23_TYPE == IRQ_TYPE_LEVEL) begin i_irq23_r <= 1'b 0;    end
      if (IRQ24_TYPE == IRQ_TYPE_LEVEL) begin i_irq24_r <= 1'b 0;    end
      if (IRQ25_TYPE == IRQ_TYPE_LEVEL) begin i_irq25_r <= 1'b 0;    end
      if (IRQ26_TYPE == IRQ_TYPE_LEVEL) begin i_irq26_r <= 1'b 0;    end
      if (IRQ27_TYPE == IRQ_TYPE_LEVEL) begin i_irq27_r <= 1'b 0;    end
      if (IRQ28_TYPE == IRQ_TYPE_LEVEL) begin i_irq28_r <= 1'b 0;    end
      if (IRQ29_TYPE == IRQ_TYPE_LEVEL) begin i_irq29_r <= 1'b 0;    end
      if (IRQ30_TYPE == IRQ_TYPE_LEVEL) begin i_irq30_r <= 1'b 0;    end
      if (IRQ31_TYPE == IRQ_TYPE_LEVEL) begin i_irq31_r <= 1'b 0;    end
      if (MEM_IRQ_TYPE == IRQ_TYPE_PULSE)
         begin
         i_irq1_r <= i_irq_a[1];    
         end
      if (INS_IRQ_TYPE == IRQ_TYPE_PULSE)
         begin
         i_irq2_r <= i_irq_a[2];    
         end
      if (IRQ3_TYPE == IRQ_TYPE_PULSE)
         begin
         if (i_swi_cancel_a[0])
           i_irq3_r <= 1'b0;
         else
           i_irq3_r <= i_irq_a[3];    
         end
      if (IRQ4_TYPE == IRQ_TYPE_PULSE)
         begin
         if (i_swi_cancel_a[1])
           i_irq4_r <= 1'b0;
         else
           i_irq4_r <= i_irq_a[4];    
         end
      if (IRQ5_TYPE == IRQ_TYPE_PULSE)
         begin
         if (i_swi_cancel_a[2])
           i_irq5_r <= 1'b0;
         else
           i_irq5_r <= i_irq_a[5];    
         end
      if (IRQ6_TYPE == IRQ_TYPE_PULSE)
         begin
         if (i_swi_cancel_a[3])
           i_irq6_r <= 1'b0;
         else
           i_irq6_r <= i_irq_a[6];    
         end
      if (IRQ7_TYPE == IRQ_TYPE_PULSE)
         begin
         if (i_swi_cancel_a[4])
           i_irq7_r <= 1'b0;
         else
           i_irq7_r <= i_irq_a[7];    
         end
      if (IRQ8_TYPE == IRQ_TYPE_PULSE)
         begin
         if (i_swi_cancel_a[5])
           i_irq8_r <= 1'b0;
         else
           i_irq8_r <= i_irq_a[8];    
         end
      if (IRQ9_TYPE == IRQ_TYPE_PULSE)
         begin
         if (i_swi_cancel_a[6])
           i_irq9_r <= 1'b0;
         else
           i_irq9_r <= i_irq_a[9];    
         end
      if (IRQ10_TYPE == IRQ_TYPE_PULSE)
         begin
         if (i_swi_cancel_a[7])
           i_irq10_r <= 1'b0;
         else
           i_irq10_r <= i_irq_a[10];  
         end
      if (IRQ11_TYPE == IRQ_TYPE_PULSE)
         begin
         if (i_swi_cancel_a[8])
           i_irq11_r <= 1'b0;
         else
           i_irq11_r <= i_irq_a[11];  
         end
      if (IRQ12_TYPE == IRQ_TYPE_PULSE)
         begin
         if (i_swi_cancel_a[9])
           i_irq12_r <= 1'b0;
         else
           i_irq12_r <= i_irq_a[12];  
         end 
      if (IRQ13_TYPE == IRQ_TYPE_PULSE)
         begin
         if (i_swi_cancel_a[10])
           i_irq13_r <= 1'b0;
         else
           i_irq13_r <= i_irq_a[13];  
         end
      if (IRQ14_TYPE == IRQ_TYPE_PULSE)
         begin
         if (i_swi_cancel_a[11])
           i_irq14_r <= 1'b0;
         else
           i_irq14_r <= i_irq_a[14];  
         end
      if (IRQ15_TYPE == IRQ_TYPE_PULSE)
         begin
         if (i_swi_cancel_a[12])
           i_irq15_r <= 1'b0;
         else
           i_irq15_r <= i_irq_a[15];  
         end
      if (IRQ16_TYPE == IRQ_TYPE_PULSE) 
         begin 
         if (i_swi_cancel_a[13])
            i_irq16_r <= 1'b0;
         else
            i_irq16_r <= i_irq_a[16];  
         end
      if (IRQ17_TYPE == IRQ_TYPE_PULSE) 
         begin 
         if (i_swi_cancel_a[14])
            i_irq17_r <= 1'b0;
         else
            i_irq17_r <= i_irq_a[17];  
         end
      if (IRQ18_TYPE == IRQ_TYPE_PULSE) 
         begin 
         if (i_swi_cancel_a[15])
            i_irq18_r <= 1'b0;
         else
            i_irq18_r <= i_irq_a[18];  
         end
      if (IRQ19_TYPE == IRQ_TYPE_PULSE) 
         begin 
         if (i_swi_cancel_a[16])
            i_irq19_r <= 1'b0;
         else
            i_irq19_r <= i_irq_a[19];  
         end
      if (IRQ20_TYPE == IRQ_TYPE_PULSE) 
         begin 
         if (i_swi_cancel_a[17])
            i_irq20_r <= 1'b0;
         else
            i_irq20_r <= i_irq_a[20];  
         end
      if (IRQ21_TYPE == IRQ_TYPE_PULSE) 
         begin 
         if (i_swi_cancel_a[18])
            i_irq21_r <= 1'b0;
         else
            i_irq21_r <= i_irq_a[21];  
         end
      if (IRQ22_TYPE == IRQ_TYPE_PULSE) 
         begin 
         if (i_swi_cancel_a[19])
            i_irq22_r <= 1'b0;
         else
            i_irq22_r <= i_irq_a[22];  
         end
      if (IRQ23_TYPE == IRQ_TYPE_PULSE) 
         begin 
         if (i_swi_cancel_a[20])
            i_irq23_r <= 1'b0;
         else
            i_irq23_r <= i_irq_a[23];  
         end
      if (IRQ24_TYPE == IRQ_TYPE_PULSE) 
         begin 
         if (i_swi_cancel_a[21])
            i_irq24_r <= 1'b0;
         else
            i_irq24_r <= i_irq_a[24];  
         end
      if (IRQ25_TYPE == IRQ_TYPE_PULSE) 
         begin 
         if (i_swi_cancel_a[22])
            i_irq25_r <= 1'b0;
         else
            i_irq25_r <= i_irq_a[25];  
         end
      if (IRQ26_TYPE == IRQ_TYPE_PULSE) 
         begin 
         if (i_swi_cancel_a[23])
            i_irq26_r <= 1'b0;
         else
            i_irq26_r <= i_irq_a[26];  
         end
      if (IRQ27_TYPE == IRQ_TYPE_PULSE) 
         begin 
         if (i_swi_cancel_a[24])
            i_irq27_r <= 1'b0;
         else
            i_irq27_r <= i_irq_a[27];  
         end
      if (IRQ28_TYPE == IRQ_TYPE_PULSE) 
         begin 
         if (i_swi_cancel_a[25])
            i_irq28_r <= 1'b0;
         else
            i_irq28_r <= i_irq_a[28];  
         end
      if (IRQ29_TYPE == IRQ_TYPE_PULSE) 
         begin 
         if (i_swi_cancel_a[26])
            i_irq29_r <= 1'b0;
         else
            i_irq29_r <= i_irq_a[29];  
         end
      if (IRQ30_TYPE == IRQ_TYPE_PULSE) 
         begin 
         if (i_swi_cancel_a[27])
            i_irq30_r <= 1'b0;
         else
            i_irq30_r <= i_irq_a[30];  
         end
      if (IRQ31_TYPE == IRQ_TYPE_PULSE) 
         begin 
         if (i_swi_cancel_a[28])
            i_irq31_r <= 1'b0;
         else
            i_irq31_r <= i_irq_a[31];  
         end

      if (( auxdc(aux_addr, AUX_IRQ_LEV) == 1'b 1 ) &
          ( aux_write == 1'b 1 ))
         begin
         i_aux_lev_r <= aux_dataw[31:3];    
         end
      else if (( auxdc(h_addr, AUX_IRQ_LEV) == 1'b 1 ) &
               ( aux_access == 1'b 1 ) & h_write == 1'b 1 )
         begin
         i_aux_lev_r <= h_dataw[31:3];  
         end
      if (( auxdc(aux_addr, AUX_IRQ_HINT) == 1'b 1 ) &
          ( aux_write == 1'b 1 ))
         begin
         i_aux_hint_r <= aux_dataw[4:0];    
         end
      else if (( auxdc(h_addr, AUX_IRQ_HINT) == 1'b 1 ) &
               ( aux_access == 1'b 1 ) & ( h_write == 1'b 1 ) )
         begin
         i_aux_hint_r <= h_dataw[4:0];  
         end
      end
   end

// Cancel software interrupts when zero is written to
// the 'hint' register.
//        
always @(
         i_aux_hint_r or
         aux_addr or
         aux_write or 
         aux_dataw
         )
   begin : cancel_hint_PROC
   
     i_swi_cancel_a = 29'b0;
   
     if ((( auxdc(aux_addr, AUX_IRQ_HINT) == 1'b 1 ) &&
          ( aux_write == 1'b 1 )) && (aux_dataw == 32'b0))
     begin
      case(i_aux_hint_r) 
        5'b 00011 : i_swi_cancel_a[0]  = 1'b1;
        5'b 00100 : i_swi_cancel_a[1]  = 1'b1;
        5'b 00101 : i_swi_cancel_a[2]  = 1'b1;
        5'b 00110 : i_swi_cancel_a[3]  = 1'b1;
        5'b 00111 : i_swi_cancel_a[4]  = 1'b1;
        5'b 01000 : i_swi_cancel_a[5]  = 1'b1; 
        5'b 01001 : i_swi_cancel_a[6]  = 1'b1;
        5'b 01010 : i_swi_cancel_a[7]  = 1'b1;
        5'b 01011 : i_swi_cancel_a[8]  = 1'b1;
        5'b 01100 : i_swi_cancel_a[9]  = 1'b1;
        5'b 01101 : i_swi_cancel_a[10] = 1'b1;
        5'b 01110 : i_swi_cancel_a[11] = 1'b1;
        5'b 01111 : i_swi_cancel_a[12] = 1'b1;
        5'b 10000 : i_swi_cancel_a[13] = 1'b1;
        5'b 10001 : i_swi_cancel_a[14] = 1'b1;
        5'b 10010 : i_swi_cancel_a[15] = 1'b1;
        5'b 10011 : i_swi_cancel_a[16] = 1'b1;
        5'b 10100 : i_swi_cancel_a[17] = 1'b1;
        5'b 10101 : i_swi_cancel_a[18] = 1'b1;
        5'b 10110 : i_swi_cancel_a[19] = 1'b1;
        5'b 10111 : i_swi_cancel_a[20] = 1'b1;
        5'b 11000 : i_swi_cancel_a[21] = 1'b1;
        5'b 11001 : i_swi_cancel_a[22] = 1'b1;
        5'b 11010 : i_swi_cancel_a[23] = 1'b1;
        5'b 11011 : i_swi_cancel_a[24] = 1'b1;
        5'b 11100 : i_swi_cancel_a[25] = 1'b1;
        5'b 11101 : i_swi_cancel_a[26] = 1'b1;
        5'b 11110 : i_swi_cancel_a[27] = 1'b1;
        5'b 11111 : i_swi_cancel_a[28] = 1'b1;      
      endcase // case(l_aux_hit)
     end
   end 

// Block out interrupts when:
//
// a. Another interrupt is already being processed (p2int/p3int)
// 
// b. The instruction in stage2 depends on the next instruction 
//    following immediately after it. (interrupt_holdoff).
// 
// c. An instruction is present in stage 2 or 3 which could 
//    disable the interrupt flags. This ensures that no 
//    interrupts can be taken between the disabling instruction
//    at the time when the appropriate interrupt flag has been
//    cleared.
// 
assign i_blockout_a = i_p2int_r | i_p2bint_r | i_p3int_r | 
                      interrupt_holdoff | flagu_block; 


// Process to show interrupt in the pipeline. The signal p123int is 
// only used with clock gating.
//
assign p123int = i_p1int_a | i_p2int_r | i_p2bint_r | i_p3int_r;

// Interrupts at stage 0
// Decide which interrupt will be processed on the next cycle. This
// part also determines the priority of interrupts.
//

//  priority subset (3) - highest
assign i_p0state3_nxt =
   ((i_irq_a[7]  & i_aux_lev_r[7])  == 1'b 1) ? S_IRQ7 : 
   ((i_irq_a[31] & i_aux_lev_r[31]) == 1'b 1) ? S_IRQ31 : 
   ((i_irq_a[30] & i_aux_lev_r[30]) == 1'b 1) ? S_IRQ30 : 
   ((i_irq_a[29] & i_aux_lev_r[29]) == 1'b 1) ? S_IRQ29 : 
   ((i_irq_a[28] & i_aux_lev_r[28]) == 1'b 1) ? S_IRQ28 : 
   ((i_irq_a[27] & i_aux_lev_r[27]) == 1'b 1) ? S_IRQ27 : 
   ((i_irq_a[26] & i_aux_lev_r[26]) == 1'b 1) ? S_IRQ26 : 
   ((i_irq_a[25] & i_aux_lev_r[25]) == 1'b 1) ? S_IRQ25 : 
   ((i_irq_a[24] & i_aux_lev_r[24]) == 1'b 1) ? S_IRQ24 : 
   ((i_irq_a[23] & i_aux_lev_r[23]) == 1'b 1) ? S_IRQ23 : 
   ((i_irq_a[22] & i_aux_lev_r[22]) == 1'b 1) ? S_IRQ22 : 
   ((i_irq_a[21] & i_aux_lev_r[21]) == 1'b 1) ? S_IRQ21 : 
   ((i_irq_a[20] & i_aux_lev_r[20]) == 1'b 1) ? S_IRQ20 : 
   ((i_irq_a[19] & i_aux_lev_r[19]) == 1'b 1) ? S_IRQ19 : 
       S_IRQ0; 

//  priority subset (2)
assign i_p0state2_nxt =
   ((i_irq_a[18] & i_aux_lev_r[18]) == 1'b 1) ? S_IRQ18 : 
   ((i_irq_a[17] & i_aux_lev_r[17]) == 1'b 1) ? S_IRQ17 : 
   ((i_irq_a[16] & i_aux_lev_r[16]) == 1'b 1) ? S_IRQ16 : 
   ((i_irq_a[15] & i_aux_lev_r[15]) == 1'b 1) ? S_IRQ15 : 
   ((i_irq_a[14] & i_aux_lev_r[14]) == 1'b 1) ? S_IRQ14 : 
   ((i_irq_a[13] & i_aux_lev_r[13]) == 1'b 1) ? S_IRQ13 : 
   ((i_irq_a[12] & i_aux_lev_r[12]) == 1'b 1) ? S_IRQ12 : 
   ((i_irq_a[11] & i_aux_lev_r[11]) == 1'b 1) ? S_IRQ11 : 
   ((i_irq_a[10] & i_aux_lev_r[10]) == 1'b 1) ? S_IRQ10 : 
   ((i_irq_a[9] & i_aux_lev_r[9]) == 1'b 1) ? S_IRQ9 : 
   ((i_irq_a[8] & i_aux_lev_r[8]) == 1'b 1) ? S_IRQ8 : 
   ((i_irq_a[7] & i_aux_lev_r[7]) == 1'b 1) ? S_IRQ7 : 
   ((i_irq_a[6] & i_aux_lev_r[6]) == 1'b 1) ? S_IRQ6 : 
   ((i_irq_a[5] & i_aux_lev_r[5]) == 1'b 1) ? S_IRQ5 : 
   ((i_irq_a[4] & i_aux_lev_r[4]) == 1'b 1) ? S_IRQ4 : 
   ((i_irq_a[3] & i_aux_lev_r[3]) == 1'b 1) ? S_IRQ3 : 
       S_IRQ0; 

//  priority subset (1)
assign i_p0state1_nxt =
   ((i_irq_a[7]  & (~i_aux_lev_r[7]))  == 1'b 1) ? S_IRQ7 : 
   ((i_irq_a[31] & (~i_aux_lev_r[31])) == 1'b 1) ? S_IRQ31 : 
   ((i_irq_a[30] & (~i_aux_lev_r[30])) == 1'b 1) ? S_IRQ30 : 
   ((i_irq_a[29] & (~i_aux_lev_r[29])) == 1'b 1) ? S_IRQ29 : 
   ((i_irq_a[28] & (~i_aux_lev_r[28])) == 1'b 1) ? S_IRQ28 : 
   ((i_irq_a[27] & (~i_aux_lev_r[27])) == 1'b 1) ? S_IRQ27 : 
   ((i_irq_a[26] & (~i_aux_lev_r[26])) == 1'b 1) ? S_IRQ26 : 
   ((i_irq_a[25] & (~i_aux_lev_r[25])) == 1'b 1) ? S_IRQ25 : 
   ((i_irq_a[24] & (~i_aux_lev_r[24])) == 1'b 1) ? S_IRQ24 : 
   ((i_irq_a[23] & (~i_aux_lev_r[23])) == 1'b 1) ? S_IRQ23 : 
   ((i_irq_a[22] & (~i_aux_lev_r[22])) == 1'b 1) ? S_IRQ22 : 
   ((i_irq_a[21] & (~i_aux_lev_r[21])) == 1'b 1) ? S_IRQ21 : 
   ((i_irq_a[20] & (~i_aux_lev_r[20])) == 1'b 1) ? S_IRQ20 : 
   ((i_irq_a[19] & (~i_aux_lev_r[19])) == 1'b 1) ? S_IRQ19 : 
       S_IRQ0; 

//  priority subset (0) - lowest
assign i_p0state0_nxt =
   ((i_irq_a[18] & (~i_aux_lev_r[18])) == 1'b 1) ? S_IRQ18 : 
   ((i_irq_a[17] & (~i_aux_lev_r[17])) == 1'b 1) ? S_IRQ17 : 
   ((i_irq_a[16] & (~i_aux_lev_r[16])) == 1'b 1) ? S_IRQ16 : 
   ((i_irq_a[15] & (~i_aux_lev_r[15])) == 1'b 1) ? S_IRQ15 : 
   ((i_irq_a[14] & (~i_aux_lev_r[14])) == 1'b 1) ? S_IRQ14 : 
   ((i_irq_a[13] & (~i_aux_lev_r[13])) == 1'b 1) ? S_IRQ13 : 
   ((i_irq_a[12] & (~i_aux_lev_r[12])) == 1'b 1) ? S_IRQ12 : 
   ((i_irq_a[11] & (~i_aux_lev_r[11])) == 1'b 1) ? S_IRQ11 : 
   ((i_irq_a[10] & (~i_aux_lev_r[10])) == 1'b 1) ? S_IRQ10 : 
   ((i_irq_a[9] & (~i_aux_lev_r[9])) == 1'b 1) ? S_IRQ9 : 
   ((i_irq_a[8] & (~i_aux_lev_r[8])) == 1'b 1) ? S_IRQ8 : 
   ((i_irq_a[7] & (~i_aux_lev_r[7])) == 1'b 1) ? S_IRQ7 : 
   ((i_irq_a[6] & (~i_aux_lev_r[6])) == 1'b 1) ? S_IRQ6 : 
   ((i_irq_a[5] & (~i_aux_lev_r[5])) == 1'b 1) ? S_IRQ5 : 
   ((i_irq_a[4] & (~i_aux_lev_r[4])) == 1'b 1) ? S_IRQ4 : 
   ((i_irq_a[3] & (~i_aux_lev_r[3])) == 1'b 1) ? S_IRQ3 : 
       S_IRQ0;
 

// Process to register the results of priority encoders from stage 0
// interrupt detection.
//
always @(posedge clk_ungated or posedge rst_a)
   begin : irq_hierarchy_PROC
   if (rst_a == 1'b 1)
      begin
      i_p0state3_r <= S_IRQ0;   
      i_p0state2_r <= S_IRQ0;   
      i_p0state1_r <= S_IRQ0;   
      i_p0state0_r <= S_IRQ0;   
      end
   else
      begin
      i_p0state3_r <= i_p0state3_nxt;   
      i_p0state2_r <= i_p0state2_nxt;   
      i_p0state1_r <= i_p0state1_nxt;   
      i_p0state0_r <= i_p0state0_nxt;   
      end
   end

// Interrupts at stage 1
// detect the highest priority interrupt from what was registered
// in stage 0 and now the associated interrupt enable is set, go to
// idle state if no interrupts
//
assign i_p1state_a = ( i_blockout_a == 1'b 1 ) ? S_IRQ0 :
                     ( i_irq_a[1]   == 1'b 1 ) ? S_IRQ1 : 
                     ( i_irq_a[2]   == 1'b 1 ) ? S_IRQ2 : 
                     ( i_p0state3_r != S_IRQ0 ) & ( e2flag_r == 1'b 1 ) ?
       i_p0state3_r : 
                     ( i_p0state2_r != S_IRQ0 ) & ( e2flag_r == 1'b 1 ) ?
       i_p0state2_r : 
                     ( i_p0state1_r != S_IRQ0 ) & ( e1flag_r == 1'b 1 ) ?
       i_p0state1_r : 
                     ( i_p0state0_r != S_IRQ0 ) & ( e1flag_r == 1'b 1 ) ?
       i_p0state0_r : 
       S_IRQ0; 

assign i_p1int_a = ( i_blockout_a == 1'b 0 ) & ((( i_p0state3_r != S_IRQ0 ) | 
                   ( i_p0state2_r != S_IRQ0 )) & ( e2flag_r == 1'b 1 ) | 
                   (( i_p0state1_r != S_IRQ0 ) | ( i_p0state0_r != S_IRQ0 )) & 
                   ( e1flag_r == 1'b 1 ) | ( instruction_error == 1'b 1 ) | 
                   ( i_irq_a[1] == 1'b 1 ) | ( i_irq_a[2] == 1'b 1 )) ?
       1'b 1 : 
       1'b 0;

assign i_p2int_nxt = ( en1 == 1'b 0 ) & ( en2 == 1'b 1 ) ?
       1'b 0 :
                     ( en1 == 1'b 1 ) ?
       i_p1int_a : 
       i_p2int_r;


// Interrupt at stage 2
// p2int is p1int passed down the pipeline when en1 = '1'.
// p1state is passed down the pipe when en1 = '1'.
//
always @(posedge clk_ungated or posedge rst_a)
   begin : irq_state2_PROC
   if (rst_a == 1'b 1)
      begin
      i_aux_lev12_r <= {2{1'b 0}};  
      i_p2state_r   <= S_IRQ0;  
      i_p2int_r     <= 1'b 0;   
      i_p2ilevel1_r <= 1'b 0;   
      end
   else
      begin
      if (( auxdc(aux_addr, AUX_IRQ_LV12) == 1'b 1 ) & ( aux_write == 1'b 1 ))
         begin
         if (aux_dataw[0] == 1'b 1)
            begin
            i_aux_lev12_r[0] <= 1'b 0;  
            end
         if (aux_dataw[1] == 1'b 1)
            begin
            i_aux_lev12_r[1] <= 1'b 0;  
            end
         end
      else if (( auxdc(h_addr, AUX_IRQ_LV12) == 1'b 1 ) &
               ( aux_access == 1'b 1 ) & ( h_write == 1'b 1 ))
         begin
         if (h_dataw[0] == 1'b 1)
            begin
            i_aux_lev12_r[0] <= 1'b 0;  
            end
         if (h_dataw[1] == 1'b 1)
            begin
            i_aux_lev12_r[1] <= 1'b 0;  
            end
         end // if (auxdc(h_addr, AUX_IRQ_LV12) == 1'b 1 &...

      if (hold_int_st2_a == 1'b0)
          i_p2int_r <= i_p2int_nxt;
      
      if (en1 == 1'b 1)
         begin
         i_p2state_r <= i_p1state_a;    

         // Detect level1 interrupts
         // This is used to generate the link register writeback at
         // stage 3, and for use in the load/store unit which needs
         // to check for pending loads to the link register.
         //
         if (
   (( i_p1state_a == S_IRQ31 ) & (~i_aux_lev_r[31]) == 1'b 1) | 
   (( i_p1state_a == S_IRQ30 ) & (~i_aux_lev_r[30]) == 1'b 1) | 
   (( i_p1state_a == S_IRQ29 ) & (~i_aux_lev_r[29]) == 1'b 1) | 
   (( i_p1state_a == S_IRQ28 ) & (~i_aux_lev_r[28]) == 1'b 1) | 
   (( i_p1state_a == S_IRQ27 ) & (~i_aux_lev_r[27]) == 1'b 1) | 
   (( i_p1state_a == S_IRQ26 ) & (~i_aux_lev_r[26]) == 1'b 1) | 
   (( i_p1state_a == S_IRQ25 ) & (~i_aux_lev_r[25]) == 1'b 1) | 
   (( i_p1state_a == S_IRQ24 ) & (~i_aux_lev_r[24]) == 1'b 1) | 
   (( i_p1state_a == S_IRQ23 ) & (~i_aux_lev_r[23]) == 1'b 1) | 
   (( i_p1state_a == S_IRQ22 ) & (~i_aux_lev_r[22]) == 1'b 1) | 
   (( i_p1state_a == S_IRQ21 ) & (~i_aux_lev_r[21]) == 1'b 1) | 
   (( i_p1state_a == S_IRQ20 ) & (~i_aux_lev_r[20]) == 1'b 1) | 
   (( i_p1state_a == S_IRQ19 ) & (~i_aux_lev_r[19]) == 1'b 1) | 
   (( i_p1state_a == S_IRQ18 ) & (~i_aux_lev_r[18]) == 1'b 1) | 
   (( i_p1state_a == S_IRQ17 ) & (~i_aux_lev_r[17]) == 1'b 1) | 
   (( i_p1state_a == S_IRQ16 ) & (~i_aux_lev_r[16]) == 1'b 1) | 
   (( i_p1state_a == S_IRQ15 ) & (~i_aux_lev_r[15]) == 1'b 1) | 
   (( i_p1state_a == S_IRQ14 ) & (~i_aux_lev_r[14]) == 1'b 1) | 
   (( i_p1state_a == S_IRQ13 ) & (~i_aux_lev_r[13]) == 1'b 1) | 
   (( i_p1state_a == S_IRQ12 ) & (~i_aux_lev_r[12]) == 1'b 1) | 
   (( i_p1state_a == S_IRQ11 ) & (~i_aux_lev_r[11]) == 1'b 1) | 
   (( i_p1state_a == S_IRQ10 ) & (~i_aux_lev_r[10]) == 1'b 1) | 
   (( i_p1state_a == S_IRQ9 ) & (~i_aux_lev_r[9]) == 1'b 1) | 
   (( i_p1state_a == S_IRQ8 ) & (~i_aux_lev_r[8]) == 1'b 1) | 
   (( i_p1state_a == S_IRQ7 ) & (~i_aux_lev_r[7]) == 1'b 1) | 
   (( i_p1state_a == S_IRQ6 ) & (~i_aux_lev_r[6]) == 1'b 1) | 
   (( i_p1state_a == S_IRQ5 ) & (~i_aux_lev_r[5]) == 1'b 1) | 
   (( i_p1state_a == S_IRQ4 ) & (~i_aux_lev_r[4]) == 1'b 1) | 
   (( i_p1state_a == S_IRQ3 ) & (~i_aux_lev_r[3]) == 1'b 1) | 
	1'b 0)
            //  level 1 interrupt
            begin
            i_p2ilevel1_r <= 1'b 1; 
            i_aux_lev12_r[0] <= 1'b 1;  
            end
         //  level 2 interrupt
         else if (i_p1state_a != S_IRQ0 )
            begin
            i_p2ilevel1_r <= 1'b 0; 
            i_aux_lev12_r[1] <= 1'b 1;  
            end
         //  no interrupt
         else
            begin
            i_p2ilevel1_r <= 1'b 0; 
            end

         end
      end
   end

 // Select the correct interrupt vector
 //
 // Select the interrupt vector address
 //
 always @(i_p2state_r)
      begin : int_vec_async_PROC
         case(i_p2state_r) 
           S_IRQ31 : i_int_vec_a = `IVECTOR_OFS31;
           S_IRQ30 : i_int_vec_a = `IVECTOR_OFS30;
           S_IRQ29 : i_int_vec_a = `IVECTOR_OFS29;
           S_IRQ28 : i_int_vec_a = `IVECTOR_OFS28;
           S_IRQ27 : i_int_vec_a = `IVECTOR_OFS27;
           S_IRQ26 : i_int_vec_a = `IVECTOR_OFS26;
           S_IRQ25 : i_int_vec_a = `IVECTOR_OFS25;
           S_IRQ24 : i_int_vec_a = `IVECTOR_OFS24;
           S_IRQ23 : i_int_vec_a = `IVECTOR_OFS23;
           S_IRQ22 : i_int_vec_a = `IVECTOR_OFS22;
           S_IRQ21 : i_int_vec_a = `IVECTOR_OFS21;
           S_IRQ20 : i_int_vec_a = `IVECTOR_OFS20;
           S_IRQ19 : i_int_vec_a = `IVECTOR_OFS19;
           S_IRQ18 : i_int_vec_a = `IVECTOR_OFS18;
           S_IRQ17 : i_int_vec_a = `IVECTOR_OFS17;
           S_IRQ16 : i_int_vec_a = `IVECTOR_OFS16;
           S_IRQ15 : i_int_vec_a = `IVECTOR_OFS15;
           S_IRQ14 : i_int_vec_a = `IVECTOR_OFS14;
           S_IRQ13 : i_int_vec_a = `IVECTOR_OFS13;
           S_IRQ12 : i_int_vec_a = `IVECTOR_OFS12;
           S_IRQ11 : i_int_vec_a = `IVECTOR_OFS11;
           S_IRQ10 : i_int_vec_a = `IVECTOR_OFS10;
           S_IRQ9 : i_int_vec_a = `IVECTOR_OFS9;
           S_IRQ8 : i_int_vec_a = `IVECTOR_OFS8;
           S_IRQ7 : i_int_vec_a = `IVECTOR_OFS7;
           S_IRQ6 : i_int_vec_a = `IVECTOR_OFS6;
           S_IRQ5 : i_int_vec_a = `IVECTOR_OFS5;
           S_IRQ4 : i_int_vec_a = `IVECTOR_OFS4;
           S_IRQ3 : i_int_vec_a = `IVECTOR_OFS3;
           S_IRQ2 : i_int_vec_a = `IVECTOR_OFS2;
           S_IRQ1 : i_int_vec_a = `IVECTOR_OFS1;
           default : i_int_vec_a = {(`INT_BASE_LSB) {1'b 0}};
         endcase // case(i_p2state_r)
      end // block: int_vec_mux

// Interrupts at stage 2B
// Generation of p2bint & p2bilev1.
// p2bint is p2int passed down the pipeline when en2 = '1'.
//
assign i_p2bint_nxt = ( en2 == 1'b 0 ) & ( en2b == 1'b 1 ) ?
       1'b 0 : 
                      ( en2 == 1'b 1 ) ? 
       i_p2int_r : 
       i_p2bint_r; 

// Move interrupt level and interrupt qualifier to stage 2B.
//
always @(posedge clk_ungated or posedge rst_a)
   begin : irq_state2b_sync_PROC
   if (rst_a == 1'b 1)
      begin
      i_p2bint_r <= 1'b 0;   
      i_p2bilevel1_r <= 1'b 0;   
      end
   else
      begin

      // Clock in newly generated stage 2B interrupt signal.
      //
      if (hold_int_st2_a)
        i_p2bint_r <= 1'b 0;
      else
        i_p2bint_r <= i_p2bint_nxt;
    
      // p2bilevl1 is set true when a level one interrupt passes
      // into stage 3. It is enabled by the pipeline enable en2.
      // (This logic does not explicitly handle pipeline tearing,
      // but as it is always qualified with p3int, then this is 
      // not a problem).
      //
      if (en2 == 1'b 1)
         begin
         i_p2bilevel1_r <= i_p2ilevel1_r;    
         end
      end
   end

// Interrupts at stage 3
// Generation of p3int & p3ilev1.
// p3int is p2bint passed down the pipeline when en2b = '1'.
//
assign i_p3int_nxt = ( en2b == 1'b 0 ) & ( en3 == 1'b 1 ) ? 
       1'b 0 : 
                     ( en2b == 1'b 1 ) ? 
       i_p2bint_r : 
       i_p3int_r; 

// Move interrupt level and interrupt qualifier to stage 3.
//
always @(posedge clk_ungated or posedge rst_a)
   begin : irq_state3_sync_PROC
   if (rst_a == 1'b 1)
      begin
      i_p3int_r <= 1'b 0;   
      i_p3ilevel1_r <= 1'b 0;   
      end
   else
      begin

      // Clock in newly generated stage 3 interrupt signal.
      //
      i_p3int_r <= i_p3int_nxt;
    
      // p3ilevl1 is set true when a level one interrupt passes
      // into stage 3. It is enabled by the pipeline enable en2.
      // (This logic does not explicitly handle pipeline tearing,
      // but as it is always qualified with p3int, then this is 
      // not a problem).
      //
      if (en2b == 1'b 1)
         begin
         i_p3ilevel1_r <= i_p2bilevel1_r;    
         end
      end
   end

//============================ Output drives =========================--
//
assign aux_hint  = i_aux_hint_r;
assign aux_lev   = i_aux_lev_r; 
assign aux_lv12  = i_aux_lev12_r;
assign int_vec   = {int_vector_base_r[PC_MSB : `INT_BASE_LSB],
                   i_int_vec_a};
assign p1int     = i_p1int_a;
assign p2bilev1  = i_p2bilevel1_r;
assign p2ilev1   = i_p2ilevel1_r;
assign p2bint    = i_p2bint_r; 
assign p2int     = i_p2int_r; 
assign p3ilev1   = i_p3ilevel1_r; 
assign p3int     = i_p3int_r; 

endmodule // module int_unit
